��V       ]�(}�}�(�name��abc��count�K�	increment�K
u}�(�name�� ��count�K�	increment�Kue.