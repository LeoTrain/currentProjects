���       ]�(}�}�(�name��abc��count�KM�	increment�Ku}�(�name�� ��count�K�	increment�Ku}�(�name��abc2��count�K$�	increment�K
ue.